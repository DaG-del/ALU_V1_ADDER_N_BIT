`timescale 1ns / 1ns

`include "incrementer/incrementer.v"
`include "comparator/comparator.v"
`include "clock/clock.v"
`include "full_adder_1_bit/full_adder.v"
`include "multiplexer/multiplexer.v"

module n_bit_adder (N2, N1, N0, )
