`timescale 1ns / 1ns

`include "comparator.v"

module comparator_tb;

reg A, B, C, D, E, F;

wire G;

comparator uut(A, B, C, D, E, F, G);

initial begin
	$dumpfile("comparator.vcd");
	$dumpvars(0, comparator_tb);
	
	A =  0;	B =  0;	C =  0;	D =  0;	E =  0;	F =  0;
	#1
	A =  0;	B =  0;	C =  0;	D =  0;	E =  0;	F =  1;
	#1
	A =  0;	B =  0;	C =  0;	D =  0;	E =  1;	F =  0;
	#1
	A =  0;	B =  0;	C =  0;	D =  0;	E =  1;	F =  1;
	#1
	A =  0;	B =  0;	C =  0;	D =  1;	E =  0;	F =  0;
	#1
	A =  0;	B =  0;	C =  0;	D =  1;	E =  0;	F =  1;
	#1
	A =  0;	B =  0;	C =  0;	D =  1;	E =  1;	F =  0;
	#1
	A =  0;	B =  0;	C =  0;	D =  1;	E =  1;	F =  1;
	#1
	A =  0;	B =  0;	C =  1;	D =  0;	E =  0;	F =  0;
	#1
	A =  0;	B =  0;	C =  1;	D =  0;	E =  0;	F =  1;
	#1
	A =  0;	B =  0;	C =  1;	D =  0;	E =  1;	F =  0;
	#1
	A =  0;	B =  0;	C =  1;	D =  0;	E =  1;	F =  1;
	#1
	A =  0;	B =  0;	C =  1;	D =  1;	E =  0;	F =  0;
	#1
	A =  0;	B =  0;	C =  1;	D =  1;	E =  0;	F =  1;
	#1
	A =  0;	B =  0;	C =  1;	D =  1;	E =  1;	F =  0;
	#1
	A =  0;	B =  0;	C =  1;	D =  1;	E =  1;	F =  1;
	#1
	A =  0;	B =  1;	C =  0;	D =  0;	E =  0;	F =  0;
	#1
	A =  0;	B =  1;	C =  0;	D =  0;	E =  0;	F =  1;
	#1
	A =  0;	B =  1;	C =  0;	D =  0;	E =  1;	F =  0;
	#1
	A =  0;	B =  1;	C =  0;	D =  0;	E =  1;	F =  1;
	#1
	A =  0;	B =  1;	C =  0;	D =  1;	E =  0;	F =  0;
	#1
	A =  0;	B =  1;	C =  0;	D =  1;	E =  0;	F =  1;
	#1
	A =  0;	B =  1;	C =  0;	D =  1;	E =  1;	F =  0;
	#1
	A =  0;	B =  1;	C =  0;	D =  1;	E =  1;	F =  1;
	#1
	A =  0;	B =  1;	C =  1;	D =  0;	E =  0;	F =  0;
	#1
	A =  0;	B =  1;	C =  1;	D =  0;	E =  0;	F =  1;
	#1
	A =  0;	B =  1;	C =  1;	D =  0;	E =  1;	F =  0;
	#1
	A =  0;	B =  1;	C =  1;	D =  0;	E =  1;	F =  1;
	#1
	A =  0;	B =  1;	C =  1;	D =  1;	E =  0;	F =  0;
	#1
	A =  0;	B =  1;	C =  1;	D =  1;	E =  0;	F =  1;
	#1
	A =  0;	B =  1;	C =  1;	D =  1;	E =  1;	F =  0;
	#1
	A =  0;	B =  1;	C =  1;	D =  1;	E =  1;	F =  1;
	#1
	A =  1;	B =  0;	C =  0;	D =  0;	E =  0;	F =  0;
	#1
	A =  1;	B =  0;	C =  0;	D =  0;	E =  0;	F =  1;
	#1
	A =  1;	B =  0;	C =  0;	D =  0;	E =  1;	F =  0;
	#1
	A =  1;	B =  0;	C =  0;	D =  0;	E =  1;	F =  1;
	#1
	A =  1;	B =  0;	C =  0;	D =  1;	E =  0;	F =  0;
	#1
	A =  1;	B =  0;	C =  0;	D =  1;	E =  0;	F =  1;
	#1
	A =  1;	B =  0;	C =  0;	D =  1;	E =  1;	F =  0;
	#1
	A =  1;	B =  0;	C =  0;	D =  1;	E =  1;	F =  1;
	#1
	A =  1;	B =  0;	C =  1;	D =  0;	E =  0;	F =  0;
	#1
	A =  1;	B =  0;	C =  1;	D =  0;	E =  0;	F =  1;
	#1
	A =  1;	B =  0;	C =  1;	D =  0;	E =  1;	F =  0;
	#1
	A =  1;	B =  0;	C =  1;	D =  0;	E =  1;	F =  1;
	#1
	A =  1;	B =  0;	C =  1;	D =  1;	E =  0;	F =  0;
	#1
	A =  1;	B =  0;	C =  1;	D =  1;	E =  0;	F =  1;
	#1
	A =  1;	B =  0;	C =  1;	D =  1;	E =  1;	F =  0;
	#1
	A =  1;	B =  0;	C =  1;	D =  1;	E =  1;	F =  1;
	#1
	A =  1;	B =  1;	C =  0;	D =  0;	E =  0;	F =  0;
	#1
	A =  1;	B =  1;	C =  0;	D =  0;	E =  0;	F =  1;
	#1
	A =  1;	B =  1;	C =  0;	D =  0;	E =  1;	F =  0;
	#1
	A =  1;	B =  1;	C =  0;	D =  0;	E =  1;	F =  1;
	#1
	A =  1;	B =  1;	C =  0;	D =  1;	E =  0;	F =  0;
	#1
	A =  1;	B =  1;	C =  0;	D =  1;	E =  0;	F =  1;
	#1
	A =  1;	B =  1;	C =  0;	D =  1;	E =  1;	F =  0;
	#1
	A =  1;	B =  1;	C =  0;	D =  1;	E =  1;	F =  1;
	#1
	A =  1;	B =  1;	C =  1;	D =  0;	E =  0;	F =  0;
	#1
	A =  1;	B =  1;	C =  1;	D =  0;	E =  0;	F =  1;
	#1
	A =  1;	B =  1;	C =  1;	D =  0;	E =  1;	F =  0;
	#1
	A =  1;	B =  1;	C =  1;	D =  0;	E =  1;	F =  1;
	#1
	A =  1;	B =  1;	C =  1;	D =  1;	E =  0;	F =  0;
	#1
	A =  1;	B =  1;	C =  1;	D =  1;	E =  0;	F =  1;
	#1
	A =  1;	B =  1;	C =  1;	D =  1;	E =  1;	F =  0;
	#1
	A =  1;	B =  1;	C =  1;	D =  1;	E =  1;	F =  1;
	#1	
	$display("test complete!");
end

endmodule
